/*************************************************************************
   Copyright 2008 Ray Salemi

   Licensed under the Apache License, Version 2.0 (the "License");
   you may not use this file except in compliance with the License.
   You may obtain a copy of the License at

       http://www.apache.org/licenses/LICENSE-2.0

   Unless required by applicable law or agreed to in writing, software
   distributed under the License is distributed on an "AS IS" BASIS,
   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
   See the License for the specific language governing permissions and
   limitations under the License.
**************************************************************************/
//
// Module tiny_cache_lib.cpubus_monitor_sm.fsm
//
// Created:
//          by - rsalemi.UNKNOWN (MAW-RSALEMI-LT)
//          at - 15:17:22 11/ 1/2006
//
// Generated by Mentor Graphics' HDL Designer(TM) 2006.1 (Build 56) Beta

module cpubus_monitor_sm( 
   clk, 
   cpu_data, 
   cpu_rd, 
   cpu_wr, 
   cpubus_address, 
   cpuwait, 
   reset, 
   active, 
   response, 
   trans
);


// Internal Declarations

input        clk;
input  [7:0] cpu_data;
input        cpu_rd;
input        cpu_wr;
input  [7:0] cpubus_address;
input        cpuwait;
input        reset;
output       active;
output       response;
output [2:0] trans;


wire clk;
wire [7:0] cpu_data;
wire cpu_rd;
wire cpu_wr;
wire [7:0] cpubus_address;
wire cpuwait;
wire monitor_reset;
wire reset;
reg active;
reg response;
reg [2:0] trans;
// Module Declarations
parameter NOTHING=0  ;
parameter READ =  1  ;
parameter WRITE  = 2  ;
parameter RESET = 3  ;
parameter CACHEHIT = 4;
parameter CACHEMISS = 5;
parameter CACHEWRITE = 6;
parameter CACHERESET = 7;

// State encoding
parameter 
          INIT_POS   = 4'd0,
          SYNC_SM    = 4'd1,
          INIT_NEG   = 4'd2,
          READ_NEG   = 4'd3,
          MISS_POS   = 4'd4,
          MISS_NEG   = 4'd5,
          MREAD_POS  = 4'd6,
          SWRITE_POS = 4'd7,
          WRITE_NEG  = 4'd8,
          MREAD_NEG  = 4'd9;

reg [3:0] current_state, next_state;
// pragma state_vector current_state

//-----------------------------------------------------------------
// Next State Block for machine csm
//-----------------------------------------------------------------
always @(
   clk or 
   cpu_rd or 
   cpu_wr or 
   cpuwait or 
   current_state or 
   reset
)
begin : next_state_block_proc
   case (current_state) 
      INIT_POS: begin
         if ( reset )
            next_state = INIT_NEG;
         else if (cpu_rd)
            next_state = READ_NEG;
         else
            next_state = INIT_NEG;
      end
      SYNC_SM: begin
         if (clk)
            next_state = INIT_POS;
         else if (~clk)
            next_state = INIT_NEG;
      end
      INIT_NEG: begin
         if ( cpu_wr )
            next_state = SWRITE_POS;
         else if ( reset )
            next_state = INIT_POS;
         else
            next_state = INIT_POS;
      end
      READ_NEG: begin
         if (~ cpuwait)
            next_state = INIT_POS;
         else if (cpuwait)
            next_state = MISS_POS;
      end
      MISS_POS: begin
         next_state = MISS_NEG;
      end
      MISS_NEG: begin
         next_state = MREAD_POS;
      end
      MREAD_POS: begin
         next_state = MREAD_NEG;
      end
      SWRITE_POS: begin
         next_state = WRITE_NEG;
      end
      WRITE_NEG: begin
         next_state = INIT_POS;
      end
      MREAD_NEG: begin
         next_state = INIT_POS;
      end
      default: 
         next_state = SYNC_SM;
   endcase
end // Next State Block

//-----------------------------------------------------------------
// Output Block for machine csm
//-----------------------------------------------------------------
always @(
   cpu_wr or 
   cpuwait or 
   current_state or 
   reset
)
begin : output_block_proc
   // Default Assignment
   active = 1;
   response = 0;
   trans = 3'b000;

   // Combined Actions
   case (current_state) 
      INIT_POS: begin
         active = 0;
      end
      SYNC_SM: begin
         active = 0;
      end
      INIT_NEG: begin
         active = 0;
         if ( cpu_wr ) begin
         end
         else if ( reset ) begin
            response = 1;
            trans = CACHERESET;
         end
      end
      READ_NEG: begin
         if (~ cpuwait) begin
             trans = CACHEHIT;
            response = 1;
         end
      end
      WRITE_NEG: begin
         response = 1;
         trans = CACHEWRITE;
      end
      MREAD_NEG: begin
         trans = CACHEMISS;
         response = 1;
      end
      default: begin
      end
   endcase
end // Output Block

//-----------------------------------------------------------------
// Clocked Block for machine csm
//-----------------------------------------------------------------
always @(
   clk or 
   negedge monitor_reset
) 
begin : clocked_block_proc
   begin
      current_state <= next_state;
   end
end // Clocked Block

endmodule // cpubus_monitor_sm
